module CPU(
	input MAIN_CLOCK,
	output [15:0] CURRENTADDRESS, REG_AC, REG_1, REG_2, REG_3, REG_AS, OUTPUT_FROM_RAM,
	output [7:0] INSTRUCTIONADDRESS, CURRENTINSTRUCTION,
	output [5:0] CMD,
	output PROCESS_DONE,
	output [15:0] DATA_OUT_RAM
	);

	
	wire PROCESS_FINISHED_FLAG,CPU_CLOCK;
	wire CPU_WRITE_EN, RAM_CLOCK;
	wire [7:0]  RAM_DATA, INSTRUCTION_ADDRESS,INSTRUCTION_DATA;
	wire [15:0] CPU_ADDRESS, CPU_DATA;
	wire [15:0] DATA_FROM_RAM;
	
	assign PROCESS_DONE = PROCESS_FINISHED_FLAG;
	assign CURRENTADDRESS = CPU_ADDRESS; // Debug
//	assign BUS_TO_RAM = RAM_DATA; // Debug
	assign INSTRUCTIONADDRESS = INSTRUCTION_ADDRESS; // Debug
	assign CURRENTINSTRUCTION = INSTRUCTION_DATA; // Debug
//	assign WEN = CPU_WRITE_EN; // Debug
	assign OUTPUT_FROM_RAM = CPU_DATA;// 
	assign DATA_OUT_RAM = DATA_FROM_RAM;

	processor Processor (
		.MAIN_CLOCK(MAIN_CLOCK),
		.PROCESS_FINISHED(PROCESS_FINISHED_FLAG),
		.DATA_FROM_RAM(DATA_FROM_RAM),
		.INSTRUCTION(INSTRUCTION_DATA),
		.CPU_CLOCK(CPU_CLOCK),
		.CPU_WRITE_EN(CPU_WRITE_EN),
		.CPU_ADDRESS(CPU_ADDRESS),
		.CPU_DATA(CPU_DATA),
		.REG_AC(REG_AC),
		.REG_1(REG_1),
		.REG_2(REG_2),
		.REG_3(REG_3),
		.REG_AS(REG_AS),
		.CMD(CMD),
//		.Z_Flag(Z_Flag),
		.INSTRUCTION_ADDRESS(INSTRUCTION_ADDRESS)
	);

	IROM_mul irom(
		.clock(CPU_CLOCK),
		.address(INSTRUCTION_ADDRESS),
		.q(INSTRUCTION_DATA)
	);

	DRAM dataram(
		.address(CPU_ADDRESS[7:0]),
		.clock(CPU_CLOCK),
		.q(DATA_FROM_RAM),
		.wren(CPU_WRITE_EN),
		.data(CPU_DATA)
	);

endmodule
