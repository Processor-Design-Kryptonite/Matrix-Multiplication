module CPU(
	input MAIN_CLOCK,
	output RAM_CLOCK,
	output PROCESS_DONE1,
	output [5:0] CMD1,
	output [15:0] REG_1_1,
	output [15:0] REG_2_1,
	output [15:0] REG_3_1, 
	output [15:0] REG_AS1, 
	output [15:0] DATA_OUT_RAM1, DATA_OUT_RAM2,
	output [15:0] REG_AC1, REG_AC2
	);

	
	wire PROCESS_FINISHED_FLAG1, PROCESS_FINISHED_FLAG2;
	wire CPU_CLOCK1, CPU_CLOCK2, DRAM_CLOCK;
	wire CPU_WRITE_EN1, CPU_WRITE_EN2;//, CPU_WRITE_EN3, CPU_WRITE_EN4;
	wire [7:0]  RAM_DATA, INSTRUCTION_DATA;
	wire [7:0]  INSTRUCTION_ADDRESS1, INSTRUCTION_ADDRESS2;//, INSTRUCTION_ADDRESS3,INSTRUCTION_ADDRESS4;
	wire [15:0] CPU_ADDRESS1, CPU_ADDRESS2;//, CPU_ADDRESS3, CPU_ADDRESS4;
	wire [15:0] CPU_DATA1, CPU_DATA2;//, CPU_DATA3, CPU_DATA4;
	wire [15:0] DATA_FROM_RAM1, DATA_FROM_RAM2;//, DATA_FROM_RAM3, DATA_FROM_RAM4;
	wire [15:0] REG_1_2;//, REG_1_3, REG_1_4; 
	wire [15:0] REG_2_2;//, REG_2_3, REG_2_4;
	wire [15:0] REG_3_2;//, REG_3_3, REG_3_4;  
	wire [15:0] REG_AS2;//, REG_AS3, REG_AS4;
	wire [5:0] CMD2;//, CMD3, CMD4;
	
	assign PROCESS_DONE1 = PROCESS_FINISHED_FLAG1;
	assign DATA_OUT_RAM1 = DATA_FROM_RAM1;
	assign DATA_OUT_RAM2 = DATA_FROM_RAM2;
//	assign DATA_OUT_RAM3 = DATA_FROM_RAM3;
//	assign DATA_OUT_RAM4 = DATA_FROM_RAM4;
	
	Clock_divider clock(
		.clock_in(MAIN_CLOCK),
		.clock_out(RAM_CLOCK)
		);

	processor core1 (
		.MAIN_CLOCK(RAM_CLOCK),
		.PROCESS_FINISHED(PROCESS_FINISHED_FLAG1),
		.DATA_FROM_RAM(DATA_FROM_RAM1),
		.INSTRUCTION(INSTRUCTION_DATA),
		.CPU_CLOCK(CPU_CLOCK1),
		.CPU_WRITE_EN(CPU_WRITE_EN1),
		.CPU_ADDRESS(CPU_ADDRESS1),
		.CPU_DATA(CPU_DATA1),
		.REG_AC(REG_AC1),
		.REG_1(REG_1_1),
		.REG_2(REG_2_1),
		.REG_3(REG_3_1),
		.REG_AS(REG_AS1),
		.CMD(CMD1),
		.INSTRUCTION_ADDRESS(INSTRUCTION_ADDRESS1)
	);
	
	processor core2 (
		.MAIN_CLOCK(RAM_CLOCK),
		.PROCESS_FINISHED(PROCESS_FINISHED_FLAG2),
		.DATA_FROM_RAM(DATA_FROM_RAM2),
		.INSTRUCTION(INSTRUCTION_DATA),
		.CPU_CLOCK(CPU_CLOCK2),
		.CPU_WRITE_EN(CPU_WRITE_EN2),
		.CPU_ADDRESS(CPU_ADDRESS2),
		.CPU_DATA(CPU_DATA2),
		.REG_AC(REG_AC2),
		.REG_1(REG_1_2),
		.REG_2(REG_2_2),
		.REG_3(REG_3_2),
		.REG_AS(REG_AS2),
		.CMD(CMD2),
		.INSTRUCTION_ADDRESS(INSTRUCTION_ADDRESS2)
	);
	
//	processor core3 (
//		.MAIN_CLOCK(RAM_CLOCK),
//		.PROCESS_FINISHED(PROCESS_FINISHED_FLAG3),
//		.DATA_FROM_RAM(DATA_FROM_RAM3),
//		.INSTRUCTION(INSTRUCTION_DATA),
//		.CPU_CLOCK(CPU_CLOCK3),
//		.CPU_WRITE_EN(CPU_WRITE_EN3),
//		.CPU_ADDRESS(CPU_ADDRESS3),
//		.CPU_DATA(CPU_DATA3),
//		.REG_AC(REG_AC3),
//		.REG_1(REG_1_3),
//		.REG_2(REG_2_3),
//		.REG_3(REG_3_3),
//		.REG_AS(REG_AS3),
//		.CMD(CMD3),
//		.INSTRUCTION_ADDRESS(INSTRUCTION_ADDRESS3)
//	);
//	
//	processor core4 (
//		.MAIN_CLOCK(RAM_CLOCK),
//		.PROCESS_FINISHED(PROCESS_FINISHED_FLAG4),
//		.DATA_FROM_RAM(DATA_FROM_RAM4),
//		.INSTRUCTION(INSTRUCTION_DATA),
//		.CPU_CLOCK(CPU_CLOCK4),
//		.CPU_WRITE_EN(CPU_WRITE_EN4),
//		.CPU_ADDRESS(CPU_ADDRESS4),
//		.CPU_DATA(CPU_DATA4),
//		.REG_AC(REG_AC4),
//		.REG_1(REG_1_4),
//		.REG_2(REG_2_4),
//		.REG_3(REG_3_4),
//		.REG_AS(REG_AS4),
//		.CMD(CMD4),
//		.INSTRUCTION_ADDRESS(INSTRUCTION_ADDRESS4)
//	);

	IROM_mul irom(
		.clock(CPU_CLOCK1),
		.address(INSTRUCTION_ADDRESS1),
		.q(INSTRUCTION_DATA)
	);

	memory_clock_generator data_clock(
		.MAIN_CLOCK(MAIN_CLOCK),
		.TICK(DRAM_CLOCK)
	);

	dataA dataram(
		//.address(CPU_ADDRESS1[7:0]),
		.address(CPU_ADDRESS1),
		.clk(DRAM_CLOCK),
		.write_en(CPU_WRITE_EN1),
		.data1(CPU_DATA1),
		.data2(CPU_DATA2),
//		.data3(CPU_DATA3),
//		.data4(CPU_DATA4),
		.q1(DATA_FROM_RAM1),
		.q2(DATA_FROM_RAM2)
//		.q3(DATA_FROM_RAM3),
//		.q4(DATA_FROM_RAM4)
	);

endmodule
